/*And gate*/

module mux16_gate (
    input wire [15:0] a0,
    input wire [15:0] a1,
    input wire [15:0] a2,
    input wire [15:0] a3,
    input wire [1:0] c,
    output reg [15:0] y
);
    

endmodule